module ClockDividerFF #(
  parameter CLK_IN_FREQ, CLK_OUT_FREQ,
  parameter integer DIVISOR = (CLK_IN_FREQ / CLK_OUT_FREQ) / 2, //Ajustado para apenas valores inteiros
  parameter TIMER_WIDTH = clog2(DIVISOR)
)(
  input clk_in,
  output reg clk_out = 0
);
`include "util.vh"

reg [TIMER_WIDTH:0] timer = 0;
always @(posedge clk_in) begin
  timer <= timer + 1;

  if (timer >= DIVISOR) begin
    clk_out <= ~clk_out;
    timer <= 0;
  end
end

endmodule